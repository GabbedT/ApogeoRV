`ifndef SCHEDULER_SV
    `define SCHEDULER_SV

module scheduler (
    input logic clk_i,
    input logic rst_n_i,
    input logic kill_instr_i,
);



endmodule : scheduler

`endif 