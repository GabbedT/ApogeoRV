`ifndef TEST_INCLUDE_SV
    `define TEST_INCLUDE_SV

// `define DECOMPRESSOR_DEBUG

// `define IDECODER_DEBUG

// `define BDECODER_DEBUG

// `define FDECODER_DEBUG

// `define WRITEBACK_DEBUG 

// `define CSR_DEBUG 

`endif