`ifndef CONFIGURATION_INCLUDE_SV
    `define CONFIGURATION_INCLUDE_SV

//====================================================================================
//      SYNTHESIS CONFIG
//====================================================================================

    /* Enable asyncronous reset */
//    `define ASYNC


//====================================================================================
//      CORE CONFIG
//====================================================================================

    /* Enable bit manipulation unit and B extension */
    `define BMU

    /* Enable or disable branch prediction */
    `define BRANCH_PREDICTOR 

    /* Total number of entries NOT bytes */

    `define BRANCH_PREDICTOR_DEPTH 1024

    `define BRANCH_TARGET_BUFFER_DEPTH 1024

    `define INSTRUCTION_BUFFER_SIZE 8

    `define STORE_BUFFER_DEPTH 8


//====================================================================================
//      MULTIPLIER CONFIG
//====================================================================================

    /* If "ASIC" is defined then the multiplier will automatically be generated 
     * with the appropriate number of pipeline stages.
     * 
     * If "FPGA" is defined then first the multiplier must be generated by the 
     * vendor tool, then the define with the stages number must be set based on
     * the IP pipeline configuration.
     * 
     * If the use of a generated IP is not possible then the file "multiplication_unit.sv" 
     * must be modified with the right module */

    /* Number of pipeline stages in the core integer multiplier, so 
     * if (MUL_PIPE_STAGES == 0) the multiplier will be combinational */
    `define MUL_PIPE_STAGES 2

`endif 