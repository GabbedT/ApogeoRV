// MIT License
//
// Copyright (c) 2021 Gabriele Tripi
// 
// Permission is hereby granted, free of charge, to any person obtaining a copy
// of this software and associated documentation files (the "Software"), to deal
// in the Software without restriction, including without limitation the rights
// to use, copy, modify, merge, publish, distribute, sublicense, and/or sell
// copies of the Software, and to permit persons to whom the Software is
// furnished to do so, subject to the following conditions:
// 
// The above copyright notice and this permission notice shall be included in all
// copies or substantial portions of the Software.
//
// THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS OR
// IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF MERCHANTABILITY,
// FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT. IN NO EVENT SHALL THE
// AUTHORS OR COPYRIGHT HOLDERS BE LIABLE FOR ANY CLAIM, DAMAGES OR OTHER
// LIABILITY, WHETHER IN AN ACTION OF CONTRACT, TORT OR OTHERWISE, ARISING FROM,
// OUT OF OR IN CONNECTION WITH THE SOFTWARE OR THE USE OR OTHER DEALINGS IN THE
// SOFTWARE.
// -----------------------------------------------------------------------------------------
// -----------------------------------------------------------------------------------------
// FILE NAME : vector_accumulator.sv
// DEPARTMENT : 
// AUTHOR : Gabriele Tripi
// AUTHOR'S EMAIL : tripi.gabriele2002@gmail.com
// -----------------------------------------------------------------------------------------
// RELEASE HISTORY
// VERSION : 1.0 
// DESCRIPTION : This module performs an 8 bit accumulation after the vector multiplication 
//               or a Q7 / Q15 saturation. For 16 bit multiplication with 32 bit addition
//               an accumulation followed by Q31 saturation is computed. 
// -----------------------------------------------------------------------------------------

`ifndef VECTOR_ACCUMULATOR_SV
    `define VECTOR_ACCUMULATOR_SV

`include "../../../../Include/Packages/vector_unit_pkg.sv"

module vector_accumulator (
    /* Registers control */
    input logic clk_i,
    input logic clk_en_i,
    input logic rst_n_i,
    
    /* Register destination used as accumulator */
    input logic [31:0] reg_accumulator_i,

    /* Result from the multiplier */
    input vmul_vector_t vmul_result_i,

    /* Specify the operation to execute */
    input vacc_uops_t operation_i,

    /* The inputs are valid */
    input logic data_valid_i,

    /* Specify how to divide the 32 bits 
     * operands and how to operate on them */
    input esize_t element_size_i,


    /* Result */
    output logic [31:0] result_o,
    output logic        data_valid_o,

    /* If the addition has overflowed */
    output logic overflow_flag_o
);


//----------------------//
//  ACCUMULATION LOGIC  //
//----------------------//

    /* Accumulator for 8 bit multiplication */
    logic [1:0][16:0] partial_8bit_accumulator;

    /* Two parallel sums */
    assign partial_8bit_accumulator[0] = vmul_result_i.vect4[0] + vmul_result_i.vect4[1];
    assign partial_8bit_accumulator[1] = vmul_result_i.vect4[2] + vmul_result_i.vect4[3];

    logic [17:0] accumulator_8bit;

    assign accumulator_8bit = partial_8bit_accumulator[0] + partial_8bit_accumulator[1];


    /* Accumulation with register destination */
    logic [31:0] reg_dest_accumulator;

    assign reg_dest_accumulator = reg_accumulator_i + accumulator_8bit;

    /* Register net */
    logic [31:0] reg_dest_accumulator_stg0;

        always_ff @(posedge clk_i) begin
            if (clk_en_i) begin
                reg_dest_accumulator_stg0 <= reg_dest_accumulator;
            end
        end


    /* Accumulator for 16 bit multiplication */
    logic [31:0] accumulator_16bit;
    logic        accumulator_sign_bit;

        always_comb begin 
            if (operation_i == FAS) begin 
                {accumulator_sign_bit, accumulator_16bit} = vmul_result_i.vect2[0] + vmul_result_i.vect2[1];
            end else begin
                {accumulator_sign_bit, accumulator_16bit} = reg_accumulator_i + vmul_result_i.vect2[0] + vmul_result_i.vect2[1];
            end
        end


//--------------------//
//  SATURATION LOGIC  //
//--------------------//

    /* Saturation logic for simple multiplication */
    vector_t    vmul_shifted, saturated_result;
    logic [3:0] sign_bit;
    logic       overflow_flag;

        always_comb begin : saturation_logic
            if (element_size_i == BIT16) begin
                {sign_bit[2], sign_bit[0]} = '0;

                /* Since the result of a multiplier has two times the operands number
                 * of bits, it needs to be shifted to be reduced */
                for (int i = 0; i < 2; ++i) begin
                    /* Do an arithmetic right shift and keep the sign bit */
                    {sign_bit[(i * 2) + 1], vmul_shifted.vect2[i]} = $signed(vmul_result_i.vect2[i]) >>> 15;
                end

                /* Check for saturation */
                for (int i = 0; i < 2; ++i) begin
                    /* If the result is positive (carry == 0) and the MSB is set, 
                     * then the number is bigger than 2^15 - 1. If the result is
                     * negative (carry == 1) and the MSB is not set, then the number
                     * is smaller than -2^15 */
                    if (sign_bit[(i * 2) + 1] ^ vmul_shifted.vect2[i][15]) begin
                        if (sign_bit[(i * 2) + 1]) begin
                            /* If the adder result is negative, set the result to 0x8000 */
                            saturated_result.vect2[i] = 16'h8000;
                        end else begin
                            /* If the adder result is positive, set the result to 0x7FFF */
                            saturated_result.vect2[i] = 16'h7FFF;
                        end

                        overflow_flag = 1'b1;
                    end else begin
                        saturated_result.vect2[i] = vmul_shifted.vect2[i];

                        overflow_flag = 1'b0;
                    end
                end
            end else if (element_size_i == BIT8) begin
                /* Since the result of a multiplier has two times the operands number
                 * of bits, it needs to be shifted to be reduced */
                for (int i = 0; i < 4; ++i) begin
                    /* Do an arithmetic right shift and keep the sign bit */
                    {sign_bit[i], vmul_shifted.vect4[i]} = $signed(vmul_shifted.vect4[i]) >>> 7;
                end

                for (int i = 0; i < 4; ++i) begin
                    /* If the result is positive (carry == 0) and the MSB is set, 
                     * then the number is bigger than 2^7 - 1. If the result is
                     * negative (carry == 1) and the MSB is not set, then the number
                     * is smaller than -2^7 */
                    if (sign_bit[i] ^ vmul_shifted.vect4[i][7]) begin
                        if (sign_bit[i]) begin
                            /* If the adder result is negative, set the result to 0x80 */
                            saturated_result.vect4[i] = 8'h80;
                        end else begin
                            /* If the adder result is positive, set the result to 0x7F */
                            saturated_result.vect4[i] = 8'h7F;
                        end

                        overflow_flag = 1'b1;
                    end else begin
                        saturated_result.vect4[i] = vmul_shifted.vect4[i];

                        overflow_flag = 1'b0;
                    end
                end
            end
        end : saturation_logic

    /* Register nets */ 
    vector_t saturated_result_stg0;
    logic    overflow_flag_stg0;

        always_ff @(posedge clk_i) begin
            if (clk_en_i) begin
                saturated_result_stg0 <= saturated_result;
                overflow_flag_stg0 <= overflow_flag;
            end
        end


    /* Saturation logic for multiplication with accumulation */
    logic [31:0] acc_sat_result;
    logic        acc_sat_overflow_flag;

        always_comb begin : accumulator_saturation_logic
            /* If the result is positive (carry == 0) and the MSB is set, 
             * then the number is bigger than 2^31 - 1. If the result is
             * negative (carry == 1) and the MSB is not set, then the number
             * is smaller than -2^31 */
            if (accumulator_sign_bit ^ accumulator_16bit[31]) begin 
                if (accumulator_sign_bit) begin
                    /* If the adder result is negative, set the result to 0x80000000 */
                    acc_sat_result = 32'h80000000;
                end else begin
                    /* If the adder result is positive, set the result to 0x7FFFFFFF */
                    acc_sat_result = 32'h7FFFFFFF;
                end

                /* Set overflow flag */
                acc_sat_overflow_flag = 1'b1;
            end else begin
                acc_sat_result = accumulator_16bit;

                acc_sat_overflow_flag = 1'b0;
            end
        end : accumulator_saturation_logic

    /* Register nets */ 
    vector_t acc_sat_result_stg0;
    logic    acc_sat_overflow_flag_stg0;

        always_ff @(posedge clk_i) begin
            if (clk_en_i) begin
                acc_sat_result_stg0 <= acc_sat_result;
                acc_sat_overflow_flag_stg0 <= acc_sat_overflow_flag;
            end
        end

//----------------//
//  OUTPUT LOGIC  //
//----------------//

    /* Register nets */
    vacc_uops_t operation_stg0;

    always_ff @(posedge clk_i) begin
        if (clk_en_i) begin
            operation_stg0 <= operation_i;
        end
    end

        always_comb begin
            /* Default values */
            result_o = '0;
            overflow_flag_o = 1'b0;

            case (operation_stg0)
                VACC: begin
                    /* Accumulation logic */
                    result_o = reg_dest_accumulator_stg0;
                    overflow_flag_o = 1'b0;
                end

                VSAT: begin
                    result_o = acc_sat_result_stg0;
                    overflow_flag_o = overflow_flag_stg0;
                end

                FAS, FAS_RD: begin
                    result_o = acc_sat_result_stg0;
                    overflow_flag_o = acc_sat_overflow_flag_stg0;
                end
            endcase
        end

    
    always_ff @(posedge clk_i `ifdef ASYNC or negedge rst_n_i `endif) begin
        if (!rst_n_i) begin
            data_valid_o <= 1'b0;
        end else begin
            data_valid_o <= data_valid_i;
        end
    end

endmodule : vector_accumulator

`endif 