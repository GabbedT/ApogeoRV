`ifndef CONTROL_STATUS_REGISTERS_SV
    `define CONTROL_STATUS_REGISTERS_SV

package control_status_registers_pkg;



endpackage : control_status_registers_pkg

import control_status_registers_pkg::*;

`endif 