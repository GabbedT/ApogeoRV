`ifndef TEST_INCLUDE_SV
    `define TEST_INCLUDE_SV

`define TEST_DESIGN

`endif